*-----------------------------------------------------------
*----------------CATALOGO DE COMPUERTAS---------------------
*-----------------------------------------------------------

*.include

*X1
*X2
*X3
*X4

*.end