*Librerias

.include 'Comp.sp'
.include 'Params.sp'


X1 A B Y vdd XORGate size = 1
*XNAND A B Y2 vdd NANDGate size = 1

.TRAN 1e-12 2e-6

.END