* Parametros para Deck

* Suggested Voltage for Technology to be used
.PARAM Vdd1=0.9			   
* Tecnologia
.PARAM Tech = 32e-9  
* Condicion fija
.PARAM UNIT_W = '2*Tech'	
.PARAM UNIT_L = Tech

