* Parametros para Deck

.PARAM Vdd1=0.9			   * Suggested Voltage for Technology to be used
.PARAM Tech = 32e-9         * Tecnologia
.PARAM UNIT_W = '2*Tech'	* Condicion fija
.PARAM UNIT_L = Tech

