*-----------------------------------------------------------
*----------------CATALOGO DE COMPUERTAS---------------------
*-----------------------------------------------------------

*.include
*.include '32nm.sp'

*X1
*X2
*X3
*X4

*.end
